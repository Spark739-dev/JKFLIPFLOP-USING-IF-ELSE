library verilog;
use verilog.vl_types.all;
entity jkflipflop_vlg_vec_tst is
end jkflipflop_vlg_vec_tst;
